include "control_register_block.sv"
include "general_purpose_reg_block.sv"
include "immediate_generator_block.sv"

